`timescale 1ns / 1ps


module bil265_proje_top(
input  clk,      // clock 
input  rst_n,    // active-low reset 
input  btnl_i,   // Left button 
input  btnu_i,   // Upper button 
input  btnr_i,   // Right button 
input  btnd_i,   // Down button 
input  rx_i,     // UART receive 
output reg tx_o      // UART transmit
    );



 
endmodule
